,.mcal_rd_vref_value (
{

    7'b0,
    7'b0,
    mcal_rd_vref_value[13:7],
    mcal_rd_vref_value[6:0]
}
)

,.iob_pin (
{

ddr4_cke[0],
ddr4_cs_n[0],
ddr4_bg[0],
ddr4_ba[1],
ddr4_ba[0],
ddr4_adr[16],
ddr4_adr[15],
ddr4_adr[14],
ddr4_adr[13],
ddr4_adr[12],
ddr4_adr[11],
ddr4_adr[10],
ddr4_adr[9],
ddr4_adr[8],
ddr4_adr[7],
ddr4_adr[6],
ddr4_adr[5],
ddr4_adr[4],
ddr4_ck_c[0],
ddr4_ck_t[0],
ddr4_adr[3],
ddr4_adr[2],
ddr4_adr[1],
ddr4_adr[0],
ddr4_nc[0],
ddr4_nc[1],
ddr4_nc[2],
ddr4_dq[15],
ddr4_dq[14],
ddr4_dq[13],
ddr4_dq[12],
ddr4_dqs_c[1],
ddr4_dqs_t[1],
ddr4_dq[11],
ddr4_dq[10],
ddr4_dq[9],
ddr4_dq[8],
ddr4_act_n,
ddr4_dm_dbi_n[1],
ddr4_nc[3],
ddr4_dq[7],
ddr4_dq[6],
ddr4_dq[5],
ddr4_dq[4],
ddr4_dqs_c[0],
ddr4_dqs_t[0],
ddr4_dq[3],
ddr4_dq[2],
ddr4_dq[1],
ddr4_dq[0],
ddr4_odt[0],
ddr4_dm_dbi_n[0]
}
)


